`ifndef __alu_vh__
`define __alu_vh__
	`define	ALU_NOP	 4'b0000
	`define	ALU_ADD	 4'b0000
	`define	ALU_SUB  4'b0001
    `define	ALU_MUL  4'b0010
	`define	ALU_AND  4'b0011
	`define	ALU_OR   4'b0100
	`define	ALU_XOR  4'b0101
    `define	ALU_EQ   4'b0110
    `define	ALU_NE   4'b0111
    `define	ALU_LT   4'b1000
    `define	ALU_GT   4'b1001
`endif //__alu_vh__
